module axi4_testbench;
    
    // Clock and reset
    logic clk;
    logic rst_n;
    
    // AXI4 Master Interface
    logic [31:0] m_axi_awaddr;
    logic [7:0]  m_axi_awlen;
    logic [2:0]  m_axi_awsize;
    logic [1:0]  m_axi_awburst;
    logic        m_axi_awvalid;
    logic        m_axi_awready;
    
    logic [31:0] m_axi_wdata;
    logic [3:0]  m_axi_wstrb;
    logic        m_axi_wlast;
    logic        m_axi_wvalid;
    logic        m_axi_wready;
    
    logic [1:0]  m_axi_bresp;
    logic        m_axi_bvalid;
    logic        m_axi_bready;
    
    logic [31:0] m_axi_araddr;
    logic [7:0]  m_axi_arlen;
    logic [2:0]  m_axi_arsize;
    logic [1:0]  m_axi_arburst;
    logic        m_axi_arvalid;
    logic        m_axi_arready;
    
    logic [31:0] m_axi_rdata;
    logic [1:0]  m_axi_rresp;
    logic        m_axi_rlast;
    logic        m_axi_rvalid;
    logic        m_axi_rready;
    
    // Coverage and assertions
    covergroup axi4_coverage @(posedge clk);
        write_burst: coverpoint m_axi_awlen {
            bins single = {0};
            bins burst_4 = {3};
            bins burst_8 = {7};
            bins burst_16 = {15};
        }
        
        read_burst: coverpoint m_axi_arlen {
            bins single = {0};
            bins burst_4 = {3};
            bins burst_8 = {7};
            bins burst_16 = {15};
        }
        
        write_response: coverpoint m_axi_bresp {
            bins okay = {2'b00};
            bins exokay = {2'b01};
            bins slverr = {2'b10};
            bins decerr = {2'b11};
        }
    endgroup
    
    axi4_coverage cov_inst = new();
    
    // Assertions
    property axi4_handshake_valid_ready(valid, ready);
        @(posedge clk) disable iff (!rst_n)
        valid && !ready |=> valid;
    endproperty
    
    assert property (axi4_handshake_valid_ready(m_axi_awvalid, m_axi_awready))
        else $error("AXI4 AW handshake violation");
    
    assert property (axi4_handshake_valid_ready(m_axi_wvalid, m_axi_wready))
        else $error("AXI4 W handshake violation");
    
    assert property (axi4_handshake_valid_ready(m_axi_arvalid, m_axi_arready))
        else $error("AXI4 AR handshake violation");
    
    // Clock generation
    always #5 clk = ~clk;
    
    // Test sequence
    initial begin
        clk = 0;
        rst_n = 0;
        
        // Initialize signals
        m_axi_awaddr = 0;
        m_axi_awlen = 0;
        m_axi_awsize = 3'b010; // 4 bytes
        m_axi_awburst = 2'b01; // INCR
        m_axi_awvalid = 0;
        
        m_axi_wdata = 0;
        m_axi_wstrb = 4'hF;
        m_axi_wlast = 0;
        m_axi_wvalid = 0;
        
        m_axi_bready = 1;
        
        m_axi_araddr = 0;
        m_axi_arlen = 0;
        m_axi_arsize = 3'b010;
        m_axi_arburst = 2'b01;
        m_axi_arvalid = 0;
        
        m_axi_rready = 1;
        
        // Reset sequence
        repeat(10) @(posedge clk);
        rst_n = 1;
        repeat(5) @(posedge clk);
        
        // Test single write
        axi4_write(32'h1000, 32'hDEADBEEF, 0);
        
        // Test burst write (4 beats)
        axi4_burst_write(32'h2000, 3, {32'h12345678, 32'h9ABCDEF0, 32'hFEDCBA98, 32'h76543210});
        
        // Test single read
        axi4_read(32'h1000, 0);
        
        // Test burst read (4 beats)
        axi4_burst_read(32'h2000, 3);
        
        // Error injection test
        axi4_write(32'hFFFF_FFFF, 32'h12345678, 0); // Invalid address
        
        repeat(100) @(posedge clk);
        
        $display("Functional Coverage: %0.2f%%", cov_inst.get_coverage());
        $finish;
    end
    
    // Write transaction task
    task axi4_write(input [31:0] addr, input [31:0] data, input [7:0] len);
        fork
            begin
                // Address channel
                m_axi_awaddr = addr;
                m_axi_awlen = len;
                m_axi_awvalid = 1;
                @(posedge clk iff m_axi_awready);
                m_axi_awvalid = 0;
            end
            begin
                // Data channel
                repeat(len + 1) begin
                    m_axi_wdata = data;
                    m_axi_wvalid = 1;
                    m_axi_wlast = (len == 0);
                    @(posedge clk iff m_axi_wready);
                    data = data + 1; // Increment for burst
                    len = len - 1;
                end
                m_axi_wvalid = 0;
                m_axi_wlast = 0;
            end
        join
        
        // Wait for response
        @(posedge clk iff m_axi_bvalid);
        $display("Write response: %0h", m_axi_bresp);
    endtask
    
    // Burst write task
    task axi4_burst_write(input [31:0] addr, input [7:0] len, input [31:0] data_array[]);
        fork
            begin
                m_axi_awaddr = addr;
                m_axi_awlen = len;
                m_axi_awvalid = 1;
                @(posedge clk iff m_axi_awready);
                m_axi_awvalid = 0;
            end
            begin
                for(int i = 0; i <= len; i++) begin
                    m_axi_wdata = data_array[i];
                    m_axi_wvalid = 1;
                    m_axi_wlast = (i == len);
                    @(posedge clk iff m_axi_wready);
                end
                m_axi_wvalid = 0;
                m_axi_wlast = 0;
            end
        join
        
        @(posedge clk iff m_axi_bvalid);
        $display("Burst write response: %0h", m_axi_bresp);
    endtask
    
    // Read transaction task
    task axi4_read(input [31:0] addr, input [7:0] len);
        m_axi_araddr = addr;
        m_axi_arlen = len;
        m_axi_arvalid = 1;
        @(posedge clk iff m_axi_arready);
        m_axi_arvalid = 0;
        
        repeat(len + 1) begin
            @(posedge clk iff m_axi_rvalid);
            $display("Read data: %0h, resp: %0h, last: %0b", 
                     m_axi_rdata, m_axi_rresp, m_axi_rlast);
        end
    endtask
    
    // Burst read task
    task axi4_burst_read(input [31:0] addr, input [7:0] len);
        m_axi_araddr = addr;
        m_axi_arlen = len;
        m_axi_arvalid = 1;
        @(posedge clk iff m_axi_arready);
        m_axi_arvalid = 0;
        
        for(int i = 0; i <= len; i++) begin
            @(posedge clk iff m_axi_rvalid);
            $display("Burst read[%0d]: %0h, resp: %0h, last: %0b", 
                     i, m_axi_rdata, m_axi_rresp, m_axi_rlast);
        end
    endtask
    
endmodule

